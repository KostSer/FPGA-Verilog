module VRAM_Green(addr, reset, clk, out);
   input clk, reset;
   input [13:0] addr;
   output [31:0] out;
//  RAMB18E1   : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB18E1_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB18E1: 18K-bit Configurable Synchronous Block RAM
   //           Artix-7
   // Xilinx HDL Language Template, version 2018.3

   // white line: D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B
   // black line: 10842108421084200421084210842108

   //10842108421084200421084210842108D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B
   //D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B10842108421084200421084210842108
   //D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6BD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B

   RAMB18E1 #(
      // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
      .SIM_COLLISION_CHECK("ALL"),
      // DOA_REG, DOB_REG: Optional output register (0 or 1)
      .DOA_REG(0),
      .DOB_REG(0),
      // INITP_00 to INITP_07: Initial contents of parity memory array
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_00 to INIT_3F: Initial contents of data memory array
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_02(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_05(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_08(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0B(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), // last white line of red
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), // last white line of green
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1A(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1D(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_20(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_23(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_24(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), // last white of blue
      .INIT_25(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B10842108421084200421084210842108),
      .INIT_26(256'h10842108421084200421084210842108D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B),
      .INIT_27(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6BD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B),
      .INIT_28(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B10842108421084200421084210842108),
      .INIT_29(256'h10842108421084200421084210842108D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B),
      .INIT_2A(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6BD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B),
      .INIT_2B(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B10842108421084200421084210842108),
      .INIT_2C(256'h10842108421084200421084210842108D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B),
      .INIT_2D(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6BD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B),
      .INIT_2E(256'hD6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B10842108421084200421084210842108),
      .INIT_2F(256'h10842108421084200421084210842108D6B5AD6B5AD6B5AFF5AD6B5AD6B5AD6B), //b8, end below all black
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_A, INIT_B: Initial values on output ports
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      // Initialization File: RAM initialization file
      .INIT_FILE("NONE"),
      // RAM Mode: "SDP" or "TDP" 
      .RAM_MODE("TDP"),
      // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      .READ_WIDTH_A(1'b1),                                                                 // 0-72
      .READ_WIDTH_B(0),                                                                 // 0-18
      .WRITE_WIDTH_A(0),                                                                // 0-18
      .WRITE_WIDTH_B(0),                                                                // 0-72
      // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      // SRVAL_A, SRVAL_B: Set/reset value for output
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      // Simulation Device: Must be set to "7SERIES" for simulation behavior
      .SIM_DEVICE("7SERIES"),
      // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   RAMB18E1_inst (
      // Port A Data: 16-bit (each) output: Port A data
      .DOADO(out),                 // 16-bit output: A port data/LSB data
      .DOPADOP(),             // 2-bit output: A port parity/LSB parity
      // Port B Data: 16-bit (each) output: Port B data
      .DOBDO(DOBDO),                 // 16-bit output: B port data/MSB data
      .DOPBDOP(),             // 2-bit output: B port parity/MSB parity
      // Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
      // when RAM_MODE="SDP")
      .ADDRARDADDR(addr),     // 14-bit input: A port address/Read address
      .CLKARDCLK(clk),         // 1-bit input: A port clock/Read clock
      .ENARDEN(1'b1),             // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(REGCEAREGCE),     // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset), // 1-bit input: A port set/reset
      .RSTREGARSTREG(RSTREGARSTREG), // 1-bit input: A port register set/reset
      .WEA(2'b0),                     // 2-bit input: A port write enable
      // Port A Data: 16-bit (each) input: Port A data
      .DIADI(DIADI),                 // 16-bit input: A port data/LSB data
      .DIPADIP(),             // 2-bit input: A port parity/LSB parity
      // Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
      // when RAM_MODE="SDP")
      .ADDRBWRADDR(ADDRBWRADDR),     // 14-bit input: B port address/Write address
      .CLKBWRCLK(clk),         // 1-bit input: B port clock/Write clock
      .ENBWREN(1'b0),             // 1-bit input: B port enable/Write enable
      .REGCEB(REGCEB),               // 1-bit input: B port register enable
      .RSTRAMB(RSTRAMB),             // 1-bit input: B port set/reset
      .RSTREGB(RSTREGB),             // 1-bit input: B port register set/reset
      .WEBWE(WEBWE),                 // 4-bit input: B port write enable/Write enable
      // Port B Data: 16-bit (each) input: Port B data
      .DIBDI(DIBDI),                 // 16-bit input: B port data/MSB data
      .DIPBDIP()              // 2-bit input: B port parity/MSB parity
   );

   // End of RAMB18E1_inst instantiation
endmodule
					
					